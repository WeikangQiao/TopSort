/**********************************************************************************
 This module is a user specified-width register
**********************************************************************************/
module qreg #(
    parameter integer N = 1
)
(
    input   logic                   i_clk   ,
    input	logic    [N-1:0]	    i_d     , 
    output	logic    [N-1:0]	    o_q
);

///////////////////////////////////////////////////////////////////////////////////
//Declarations
///////////////////////////////////////////////////////////////////////////////////
logic   [N-1:0]	    q_reg;

///////////////////////////////////////////////////////////////////////////////////
//Main body of the code
///////////////////////////////////////////////////////////////////////////////////
always_ff @(posedge i_clk) begin
		q_reg <= i_d;
end

assign o_q = q_reg;

endmodule