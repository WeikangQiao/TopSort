//`define USE_VIVADO_SYNTHESIS

/***** parameters                                                                     *****/
/******************************************************************************************/
/*
`define  DATA_WIDTH   (32)
`define  KEY_WIDTH    (32) 
`define  BUNDLE_WIDTH (16)
`define  INV_BUNDLE   (0) 
*/

/******************************************************************************************/
`define LOG2(x) ((x<=1)?0:\
(x<=2)?1:\
(x<=4)?2:\
(x<=8)?3:\
(x<=16)?4:\
(x<=32)?5:\
(x<=64)?6:\
(x<=128)?7:\
(x<=256)?8:\
(x<=512)?9:\
(x<=1024)?10:64)